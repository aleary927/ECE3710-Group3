/*
* Testbench for verifying RF (register file) module.
*/

module tb_RF();

  reg clk;

  reg [3:0] addr1, addr2; // addresses
  reg wr_en;        // write enable
  reg [15:0] wr_data;    // write data
  wire [15:0] rd_data1, rd_data2; // read data

  RF rf(
    .clk(clk), 
    .wr_en(wr_en), 
    .wr_data(wr_data), 
    .addr1(addr1), .addr2(addr2), 
    .rd_data1(rd_data1), .rd_data2(rd_data2));
  

  // generate clock signal
  initial begin
    clk = 0;
    forever #5 clk = ~clk;
  end

  // instanciate inputs
  initial begin
    addr1 = 0;
    addr2 = 0;
    wr_data = 0;
    wr_en = 0;
  end

  // main testbench code
  initial begin
    $display("Starting testbench for RF (register file)");

    // ===================
    // TEST WRITING TO RF
    // ===================

    // test simple write
    addr1 = 5;
    wr_en = 1;
    wr_data = 1000;
    #10;
    if (rf.registers[addr1] != wr_data)
      $display("error: result not written to register when write enabled");

    // test not writing when write enable not high
    addr1 = 6;
    wr_en = 0;
    #10;
    if (rf.registers[addr1] == wr_data)
      $display("error: unexpected write to register when write not enabled");

    // perform write so that there is data for further tests
    wr_en = 1;
    wr_data = 45;
    #10;
    wr_en = 0;

    // =========================
    // TEST READING FROM RF
    // =========================

    // test reading from 2 different registers
    addr1 = 5;
    addr2 = 6;
    #10;
    if (rd_data1 != rf.registers[addr1] || rd_data2 != rf.registers[addr2])
      $display("error: dual read did not function properly");

    // test reading from same register
    addr2 = addr1;
    #10;
    if (rd_data1 != rf.registers[addr1] || rd_data2 != rf.registers[addr1])
      $display("error: reading from same address did not function properly");

    
    $display("testbench complete");
  end

endmodule
