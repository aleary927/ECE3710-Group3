/*
* Control FSM for CR16 CPU.
*/
module CPU_Controller(); 

endmodule
