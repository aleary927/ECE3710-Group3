module VGA (input clk, 
				output [7:0]VGA_RED, VGA_GREEN, VGA_BLUE, 
				output VGA_CLK,     // VGA pixel clock (25MHz)
				output VGA_BLANK_N, // Active-low blanking signal
				output VGA_HS,      // Horizontal sync output
				output VGA_SYNC_N, // assign low
				output VGA_VS);       // added here for desired T-Bird behavior

	// here will be using h_count and v_count and bright for pixels 
	// connect hsync and vsync to VGA_HS and VGA_VS signals 

	 wire hSync, vSync, bright;
    wire [9:0] hCount, vCount;
	 wire En; 
	 
	 wire [2:0] rgb; 
	 
	 reg [3:0] new_tile = 4'b0000; 
	 
	 
	  reg rst = 0; 
	 
	 
	 wire[3:0] dead; 
	 
	 
	 
	 
	 // CODE TO GENERATE TILES ON A REGULAR BASIS

    parameter MAX_COUNT = 100000000; // 250,000,000 cycles

    reg [27:0] counter; // 28-bit counter to count clock cycles

    always @(posedge clk) begin
		rst = 0;
    if (counter >= MAX_COUNT - 1) begin
        counter <= 0; // Reset counter
        // Update new_tile signal to generate new tile
        if (new_tile == 4'b0000)
            new_tile <= 4'b0001;
        else if (new_tile == 4'b0001)
            new_tile <= 4'b0011;
        else if (new_tile == 4'b0011)
            new_tile <= 4'b0111;
        else if (new_tile == 4'b0111)
            new_tile <= 4'b1111;
        else
            new_tile <= 4'b0001; // Reset new_tile
        rst = 1;
		end else begin
        counter <= counter + 1; // Increment counter
		end
	end
	 
	 
	 
	 
	 
	 parameter NUM_LANES = 4;       // Number of lanes
  //  parameter MAX_TILES = 10;      // Maximum number of tiles per lane
	 
	 // TRACK ALL TILES position
	                           // 4 lanes     // 10 tiles max per lane
	// wire [9:0] y_pos [NUM_LANES-1:0];//[MAX_TILES-1:0];
	 
	wire [9:0] y_pos_one; 
	wire [9:0] y_pos_two; 
	wire [9:0] y_pos_three; 
	wire [9:0] y_pos_four; 
	 
	 
	SlowMover mover_one (
	 .clk(clk), 
	 .live(new_tile[0]),
    .y_pos(y_pos_one), 
	// .dead(dead[0])
	);
	
	SlowMover mover_two (
	 .clk(clk), 
	 .live(new_tile[1]),
    .y_pos(y_pos_two), 
	// .dead(dead[1])
	);
	
	SlowMover mover_three (
	 .clk(clk), 
	 .live(new_tile[2]),	 
    .y_pos(y_pos_three), 
	 //.dead(dead[2])
	);
	
	SlowMover mover_four (
	 .clk(clk),   
	 .live(new_tile[3]),	 
    .y_pos(y_pos_four), 
	// .dead(dead[3])
	);
	


	 
	 
	 
	 

    // Instantiate the vgaControl module
    vgaControl vgaInst (
        .clk(clk),       
        .clr(1'b1),       
        .hSync(hSync),   
        .vSync(vSync),    
        .bright(bright),  
        .hCount(hCount),   
        .vCount(vCount),   
		  .En(En)       //vga clock
    );
		 
		 
		 // Instantiate the bitGen_Glyph module
	bitGen_Glyph glyph_inst (
		 .clk(clk),                 
		 .live_tile(new_tile),     
		 .h_count(hCount),           
		 .v_count(vCount), 
		 .y_pos_one(y_pos_one),
		 .y_pos_two(y_pos_two),
		 .y_pos_three(y_pos_three),
		 .y_pos_four(y_pos_four),
		 .rgb(rgb)                   
	);
	

	 
	 

	 
	 assign VGA_CLK = En;        // My 25Mhz clock
											 
	 assign VGA_SYNC_N = 1'b0;
	 
    assign VGA_BLANK_N = bright; // Active low signal: invert the bright signal for blanking
    assign VGA_HS = hSync;       // Connect horizontal sync
    assign VGA_VS = vSync;       // Connect vertical sync
	 
	 
	 assign VGA_RED = {8{rgb[2]}}; // concatenate each to 8 bit value. 
	 assign VGA_GREEN = {8{rgb[1]}}; 
	 assign VGA_BLUE = {8{rgb[0]}}; 


endmodule



	
module bitGen_Glyph (
    input clk,                // System clock
	 input [3:0] live_tile, 
    input [9:0] h_count,      // Current pixel x-coordinate
    input [9:0] v_count,      // Current pixel y-coordinate
	 input [9:0] y_pos_one, //[NUM_LANES-1:0], //[MAX_TILES-1:0]
	 input [9:0] y_pos_two,
	 input [9:0] y_pos_three,
	 input [9:0] y_pos_four,
    output reg [2:0] rgb      // RGB output
);

    // Parameters for screen and lane dimensions
    parameter SCREEN_WIDTH = 640;
    parameter SCREEN_HEIGHT = 480;
    parameter NUM_LANES = 6;                     // Number of black lanes
    parameter LANE_WIDTH = SCREEN_WIDTH / NUM_LANES; // Width of each lane
    parameter LINE_WIDTH = 2;                   // Thickness of the white lines
	 
	 parameter BLOCK_LENGTH = 90; 
	 
	 
		//reg [9:0] beg_y_pos; 
	   wire [9:0] y_position;
		
		//wire [3:0] live_lane; 

    // Instantiate SlowMover to generate the Y position for the block
//    SlowMover slow_mover_inst (
//        .clk(clk),          // Connect the system clock
//        .y_pos(y_position)  // Receive the Y-coordinate
//    );
//	 
	 

    always @(*) begin
        // Default background color: black
        rgb = 3'b000; // Black
		  
		  if(h_count <(106)) begin 
					rgb = 3'b011;
		  end 
		  
		  
		  if((h_count >= 106 && h_count < 108) ||
			 (h_count >= 212 && h_count < 214) ||
			 (h_count >= 318 && h_count < 320) ||
			 (h_count >= 424 && h_count < 426) ||
			 (h_count >= 528 && h_count < 530)) begin
			 rgb = 3'b111; // White
		  end
		  

		  if (h_count >= 108 && h_count < 212 && v_count >= 450) begin
				 rgb = 3'b100;
			end
			else if (h_count >= 214 && h_count < 318 && v_count >= 450) begin
				 rgb = 3'b101;
			end
			else if (h_count >= 320 && h_count < 424 && v_count >= 450) begin
				 rgb = 3'b010;
			end
			else if (h_count >= 426 && h_count < 528 && v_count >= 450) begin
				 rgb = 3'b110;
			end

		  
		  if(h_count >= (530)) begin 
					rgb = 3'b011;
		  end 
		  
		  
		
		// loop y_position[0]
    if (live_tile[0] && h_count >= 108 && h_count < 212 && 
        v_count >= y_pos_one && v_count < y_pos_one + BLOCK_LENGTH && (y_pos_one + BLOCK_LENGTH) < 450) begin
		  
		  
        rgb = 3'b111; 
    end

		 // loop y_position [1]
    if (live_tile[1] && h_count >= 214 && h_count < 318 && 
        v_count >= y_pos_two && v_count < y_pos_two + BLOCK_LENGTH && (y_pos_two + BLOCK_LENGTH) < 450) begin
        rgb = 3'b111; 
    end

  
		// loop y_position [2]
    if (live_tile[2] && h_count >= 320 && h_count < 424 && 
        v_count >= y_pos_three && v_count < y_pos_three + BLOCK_LENGTH && (y_pos_three + BLOCK_LENGTH) < 450) begin
        rgb = 3'b111; 
    end

 
	 // loop y_position [3]
    if (live_tile[3] && h_count >= 426 && h_count < 528 && 
        v_count >= y_pos_four && v_count < y_pos_four + BLOCK_LENGTH && (y_pos_four + BLOCK_LENGTH) < 450) begin
        rgb = 3'b111; 

end

		  
		  
		  
      
    end

endmodule

















module SlowMover(
    input clk,               
    input live,               
    output reg [9:0] y_pos    // Y-coordinate of the block
);

    parameter BLOCK_LENGTH = 90; 
    parameter CLOCK_FREQ = 50000000;     
    parameter BLOCK_SPEED = 70;            // 70 pixels/second
    parameter MAX_COUNT = CLOCK_FREQ / BLOCK_SPEED; // Cycles per Y increment

    reg [25:0] counter; // 26-bit counter for clock cycles

    // Initialize signals
    initial begin
        y_pos = 0;
        counter = 0;
    end

    always @(posedge clk) begin
        if (!live) begin
            // If not live, reset counters
            counter <= 0;
        end else begin
            // Increment counter and update Y-position
            if (counter >= MAX_COUNT - 1) begin
                counter <= 0;           // Reset counter
                y_pos <= y_pos + 1;     // Increment Y-position
            end else begin
                counter <= counter + 1; // Increment counter
            end

            // Reset Y-position if the block goes out of bounds
            if ((y_pos + BLOCK_LENGTH) > 450) begin
                y_pos <= 0; // Reset to top
            end
        end
    end

endmodule



































//
//
////BLOCK LOGIC MODULE
//module SlowMover(
//    input clk,                // 50 MHz clock
//	 input rst,  
//	 input [3:0] new_tile,
//	 output reg [3:0] live_tile, 
//    output reg [9:0] y_pos [3:0]//[MAX_TILES-1:0] // 2D array for Y-coordinates of tiles
//);
//
//    // Parameters
//    parameter NUM_LANES = 4;       // Number of lanes
//   // parameter MAX_TILES = 10;      // Maximum number of tiles per lane
//    parameter BLOCK_LENGTH = 90;   // Length of each block
//    parameter SCREEN_HEIGHT = 480; // Height of the screen
//    parameter CLOCK_FREQ = 50_000_000;      // 50 MHz clock
//    parameter BLOCK_SPEED = 50;             // 50 pixels/second
//    parameter MAX_COUNT = CLOCK_FREQ / BLOCK_SPEED; // Cycles per Y increment
//
//    // 2D array for counters
//    reg [25:0] counter [NUM_LANES-1:0]; ///[MAX_TILES-1:0];
//	 
//
//    // Initialize arrays
//    integer lane; 
//	
//	 
//
//    // Always block to update positions
//    always @(posedge clk ) begin
//	 
//		if(rst) live_tile <= 4'b0000; 
//	 
//	 
//	   else begin
//	 
//        for (lane = 0; lane < NUM_LANES; lane = lane + 1) begin
//			   if(new_tile[lane] == 1) begin
//				
//					//live_tile[lane] <= 1; 
//				 
//                if (counter[lane] >= MAX_COUNT - 1) begin
//                    counter[lane] <= 0; // Reset counter
//                    y_pos[lane] <= y_pos[lane] + 1; // Increment Y-position
//                end else begin
//                    counter[lane] <= counter[lane] + 1; // Increment counter
//                end
//
//                // Make block disappear if it exceeds screen height for now got ot hte top
//                if ((y_pos[lane] + BLOCK_LENGTH) > SCREEN_HEIGHT) begin
//							y_pos[lane] <= 0; 
//							//live_tile[lane] <= 0; 
//                end
//				  end 
//				  
//				  
//				  //else live_tile[lane] <= 0; 
//			end
//		  
//		  end
//    end
//
//endmodule







