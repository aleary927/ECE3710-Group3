module ALU #(parameter DATA_WIDTH)
  (
  input [DATA_WIDTH - 1:0] a,
  input [DATA_WIDTH - 1:0] b,
  input [2:0] select,
  output [DATA_WIDTH - 1:0] out,
  output C, L, F, Z, N
  );


endmodule
