/* 
* Highest level file. 
* This file links the CPU and all external components (I/O and memory).
*/
module System(
  input clk,
  input reset,

  // vga outputs

  // other I/O outputs / inputs
); 

  // CPU 
  // I/O mapped memory 
  // VGA controller

endmodule
